	* BJT SCHMITT TRIGGER

	VDD		1 0		5V
	VIN		4 0		PULSE (0V 5V 0S 0.5US 0.5US 0S 1.0US)

	R1		1 2		2K
	R2		1 3		1.2K
	R3		5 0		460

	Q1		2 4 5	Q2N3904
	Q2		3 2 5	Q2N3904

	*		Model for 2N3904 NPN BJT (from Eval library in Pspice)
	.model Q2N3904	NPN(Is=6.734f Xti=3 Eg=1.11 Vaf=74.03 Bf=416.4 Ne=1.259
	+		Ise=6.734f Ikf=66.78m Xtb=1.5 Br=.7371 Nc=2 Isc=0 Ikr=0 Rc=1
	+		Cjc=3.638p Mjc=.3085 Vjc=.75 Fc=.5 Cje=4.493p Mje=.2593 Vje=.75
	+		Tr=239.5n Tf=301.2p Itf=.4 Vtf=4 Xtf=2 Rb=10)

	.TRAN	0.1US 2.0US

	.PROBE
	.END
