* DOUBLE BUFFERED 2-INPUT NOR GATE

VDD		2 0			5V
VIN		5 0			PULSE (0 5 0 0.001NS 0.001NS 0.10MS 0.24MS)

MP1		6 5 2 2		PMOD1
MP2		4 5 6 2		PMOD1
MP3		3 4 2 2		PMOD2
MP4		1 3 2 2		PMOD3

MN1		4 5 0 0		NMOD1
MN2		4 5 0 0		NMOD1
MN3		3 4 0 0		NMOD2
MN4		1 3 0 0		NMOD3

C		1 0			0.1UF

*** NMOS MODELS ***

.MODEL NMOD1 NMOS (L=5U W=10U KP=69U GAMMA=0.37
+LAMBDA=0.06 RD=1 RS=1 VTO=1.0 TOX=0.04U
+CBD=2F CBS=2F CJ=200U CGBO=200P CGSO=40P CGDO=40P)

.MODEL NMOD2 NMOS (L=5U W=40U KP=69U GAMMA=0.37
+LAMBDA=0.06 RD=1 RS=1 VTO=1.0 TOX=0.04U
+CBD=2F CBS=2F CJ=200U CGBO=200P CGSO=40P CGDO=40P)

.MODEL NMOD3 NMOS (L=5U W=100U KP=69U GAMMA=0.37
+LAMBDA=0.06 RD=1 RS=1 VTO=1.0 TOX=0.04U
+CBD=2F CBS=2F CJ=200U CGBO=200P CGSO=40P CGDO=40P)

*** PMOS MODELS ***

.MODEL PMOD1 PMOS (L=5U W=50U KP=34.5U GAMMA=-0.37
+LAMBDA=0.06 RD=1 RS=1 VTO=-1.0 TOX=0.04U
+CBD=2F CBS=2F CJ=200U CGBO=200P CGSO=40P CGDO=40P)

.MODEL PMOD2 PMOS (L=5U W=100U KP=34.5U GAMMA=-0.37
+LAMBDA=0.06 RD=1 RS=1 VTO=-1.0 TOX=0.04U
+CBD=2F CBS=2F CJ=200U CGBO=200P CGSO=40P CGDO=40P)

.MODEL PMOD3 PMOS (L=5U W=250U KP=34.5U GAMMA=-0.37
+LAMBDA=0.06 RD=1 RS=1 VTO=-1.0 TOX=0.04U
+CBD=2F CBS=2F CJ=200U CGBO=200P CGSO=40P CGDO=40P)

.TRAN	0.001MS 0.48MS

.PROBE
.END