* CMOS INVERTER
VDD 1 0 10
VIN 2 0

MP 3 2 1 1 PE
MN 3 2 0 0 NE

.MODEL PE PMOS (VTO=-2.7 KP=380E-6)
.MODEL NE NMOS (VTO=3.0 KP=560E-6)
.DC VIN 0 10 0.05
.PROBE
.END
