* DELAY FLIP-FLOP

.include "C:\Program Files\OrCAD\OrCAD_16.6_Lite\tools\pspice\library\dig_io.lib"
.include "C:\Program Files\OrCAD\OrCAD_16.6_Lite\tools\pspice\library\7400.lib"

VCLK	1 0		PULSE (0.5V 2.5V 0S 0.1NS 0.1NS 2MS 4MS)
VD		2 0		PULSE (0.5V 2.5V 0.1MS 0.1NS 0.1NS 5MS 10MS)

X1		2 1 3	7400
X2		1 3 4	7400
X3		3 6 5	7400
X4		4 5 6	7400

R1		5 0		10K
R2		6 0		10K

.TRAN	0.001MS 50MS
.PROBE
.END
