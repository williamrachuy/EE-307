* PMOS CURRENT VS. VOLTAGE CHARACTERISTICS
VSD 1 0
VGS 2 0
MP 0 2 1 0 PE

.MODEL PE PMOS (VTO=-2.7 KP=380E-6)
.DC VSD 0 -10 0.05 VGS 0 -10 2
.PROBE
.END