* P7.2 RD = 100K

VDD 1 0 5
VIN	2 0
RD	1 3 100K
MD	3 2 0 0 NMOD1

.MODEL NMOD1 NMOS (KP=200E-6 VTO=1.0)

.DC VIN 0 5 10m

.PROBE
.END
