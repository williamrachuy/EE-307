* EXPERIMENT 2 PRELAB SIMULATION: FIGURE 2.2b
VDD 1 0 5
VIN 2 0
RL  1 4 5.1K
ML  4 4 3 0 NMOD1
MD  3 2 0 0 NMOD1

.MODEL NMOD1 NMOS (L=3U W=6U KP=69U GAMMA=0.37
+LAMBDA=0.06 RD=1 RS=1 VTO=1.0 TOX=0.04U
+CBD=2F CBS=2F CJ=200U CGBO=200P CGSO=40P CGDO=40P)

.MODEL PMOD1 PMOS (L=3U W=6U KP=34.5U GAMMA=-0.37
+LAMBDA=0.06 RD=1 RS=1 VTO=-1.0 TOX=0.04U
+CBD=2F CBS=2F CJ=200U CGBO=200P CGSO=40P CGDO=40P)

.DC VIN 0 5 0.05

.PROBE
.END