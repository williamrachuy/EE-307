* NMOS CURRENT VS. VOLTAGE CHARACTERISTICS
VDS 1 0
VGS 3 0
MN 1 3 0 0 NE

.MODEL NE NMOS (VTO=3 KP=560E-6)
.DC VDS 0 20 0.05 VGS 0 10 2
.PROBE
.END
