* ONE-STAGE OF A DYNAMIC CMOS SHIFT REGISTER

VDD		8 0			5

V1		6 0			PULSE (5 0 0 0.1NS 0.1NS 2MS 4MS)
V2		7 0			PULSE (0 5 1MS 0.1NS 0.1NS 2MS 4MS)
VIN		4 0			PULSE (0 5 0 0.1NS 0.1NS 8MS 16MS)

MP1		5 1 8 8		PMOD1
MP2		3 2 8 8		PMOD1
MP3		4 3 8 8		PMOD1
MP4		4 6 1 1		PMOD1
MP5		5 7 2 2		PMOD1

MN1		5 1 0 0		NMOD1
MN2		3 2 0 0		NMOD1
MN3		4 3 0 0		NMOD1
MN4		4 7 1 1		NMOD1
MN5		5 6 2 2		NMOD1

.MODEL PMOD1 PMOS (L=3U W=6U KP=34.5U GAMMA=-0.37
+LAMBDA=0.06 RD=1 RS=1 VTO=-1.0 TOX=0.04U
+CBD=2F CBS=2F CJ=200U CGBO=200P CGSO=40P CGDO=40P)

.MODEL NMOD1 NMOS (L=3U W=6U KP=69U GAMMA=0.37
+LAMBDA=0.06 RD=1 RS=1 VTO=1.0 TOX=0.04U
+CBD=2F CBS=2F CJ=200U CGBO=200P CGSO=40P CGDO=40P)

.TRAN 0.001MS 16MS

.PROBE
.END