* 6.2a
VDD  1 0 5
VI 3 0 4
ML 1 1 2 2 NEL
MD 2 3 0 0 NED

.MODEL NEL NMOS (VTO=1 KP=100E-6)
.MODEL NED NMOS (VTO=1 KP=200E-6)
.END