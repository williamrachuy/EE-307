* FIG 7.8

MP1		3 2 1 1 PCH
MP2		5 4 3 1 PCH
MN1		5 2 0 0 NCH
MN2		5 4 0 0 NCH

VA		2 0
VB		4 0 0
VDD		1 0 DC 5

.PROBE
.MODEL PCH PMOS (VTO = -1.0 KP = 25E-6 GAMMA = 0.4)
.MODEL NCH NMOS (VTO = 1.0 KP = 50E-6 GAMMA = 0.4)
.DC VA 0 5V 0.1V
.END
