* P7.3

VDD 1 0 5
VIN	4 0
ML	1 1 3 3 NMODL
MD	3 4 0 0 NMODD

.MODEL NMODL NMOS (KP=20E-6 VTO=1.0)
.MODEL NMODD NMOS (KP=100E-6 VTO=1.0)

.DC VIN 0 5 10m

.PROBE
.END
