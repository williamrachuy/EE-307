* P7.11

VDD 1 0 10
VIN	2 0
MP	3 2 1 1 PMOD
MN	3 2 0 0 NMOD

.MODEL PMOD PMOS (KP=20E-6 VTO=-1.0)
.MODEL NMOD NMOS (KP=80E-6 VTO=0.8)

.DC VIN 0 10 10m

.PROBE
.END
