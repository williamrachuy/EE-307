* TTL INVERTER WITH CAPACITIVE LOAD

VDD		1 0		5
VIN		2 0		PULSE (0 5 0 1NS 1NS 0.5MS 1MS)

R1		1 5		1.5K
R2		9 0		1.0K
RB		1 4		3.9K
RC		1 6		0.1K

Q1		7 4 2	BJTMOD
Q2		5 7 9	BJTMOD
Q3		3 9 0	BJTMOD
Q4		6 5 8	BJTMOD

D1		8 3		D1

C		3 0		20P

.MODEL BJTMOD NPN (BF=156 BR=0.1 VAF=100 VAR=100
+VJC=0.75 VJE=0.75 TF=0.28P TR=10N CJE=1.02P CJC=0.99P)

.MODEL D1 D RS=1 IS=1E-15

.TRAN 0.1US 100MS

.PROBE
.END