* CMOS INVERTER WITH CAPACITIVE LOAD

VDD		1 0			5
VIN		2 0			PULSE (0 5 0 1NS 1NS 1.5MS 4MS)
MP		3 2 1 1		PMOD
MN		3 2 0 0 	NMOD
C		3 0			0.1UF

.MODEL NMOD NMOS (L=3U W=6U KP=69U GAMMA=0.37
+LAMBDA=0.06 RD=1 RS=1 VTO=1.0 TOX=0.04U
+CBD=2F CBS=2F CJ=200U CGBO=200P CGSO=40P CGDO=40P)

.MODEL PMOD PMOS (L=3U W=6U KP=34.5U GAMMA=-0.37
+LAMBDA=0.06 RD=1 RS=1 VTO=-1.0 TOX=0.04U
+CBD=2F CBS=2F CJ=200U CGBO=200P CGSO=40P CGDO=40P)

.TRAN	0.1MS 12MS 4MS

.PROBE
.END