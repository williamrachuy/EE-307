* BICMOS INVERTER WITH CAPACITIVE LOAD

VDD		1 0			5V
VIN		6 0			PULSE (0 5 0 1NS 1NS 20US 40US)

QMOS6	3 2 1 1		PMOD
QMOS3	0 2 3 3		PMOD
QMOS4	4 2 5 5		NMOD
QMOS2	5 3 0 0		NMOD

QBJT4	1 3 4		BJTMOD
QBJT5	4 5 0		BJTMOD

CL		4 0			0.1UF

.MODEL NMOD NMOS (L=3U W=6U KP=69U GAMMA=0.37
+LAMBDA=0.06 RD=1 RS=1 VTO=1.0 TOX=0.04U
+CBD=2F CBS=2F CJ=200U CGBO=200P CGSO=40P CGDO=40P)

.MODEL BJTMOD NPN (BF=156 BR=0.1 VAF=100 VAR=100
+VJC=0.75 VJE=0.75 TF=0.28P TR=10N CJE=1.02P CJC=0.99P)

.TRAN	0.1US 80US

.PROBE
.END
